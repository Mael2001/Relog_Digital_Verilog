module Controlador_MILSEG(
    input [6:0] MILSEG,
    input CLK,
    input ALARM,
    //Digito Izquierda
    output reg A7,
    output reg B7,
    output reg C7,
    output reg D7,
    output reg E7,
    output reg F7,
    output reg G7,
    output reg DP7,
    //Digito Derecho
    output reg A8,
    output reg B8,
    output reg C8,
    output reg D8,
    output reg E8,
    output reg F8,
    output reg G8,
    output reg DP8
);
initial begin
    //Izquierda
    A7=0;
    B7=0;
    C7=0;
    D7=0;
    E7=0;
    F7=0;
    G7=0;
    DP7=0;
    //Derecha
    A8=0;
    B8=0;
    C8=0;
    D8=0;
    E8=0;
    F8=0;
    G8=0;
    DP8=0;
end

    reg[5:0] numero;

always @(posedge CLK)
begin
    if(ALARM)
    begin
        numero<=0;
    end
    else
    begin
        numero<=MILSEG;
    end
 case(numero)
 0:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 1:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 2:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 3:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 4:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 5:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 6:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 7:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 8:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 9:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 10:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 11:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 12:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 13:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 14:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 15:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 16:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 17:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 18:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 19:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 20:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 21:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 22:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 23:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 24:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;  
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 25:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;  
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 26:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;  
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 27:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;  
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;   
 end
 28:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1;  
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 29:
 begin
     
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=0;
    D7<=1;
    E7<=1;
    F7<=0;
    G7<=1; 
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1; 
 end
 30:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 31:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 32:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 33:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;   
 end
 34:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 35:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 36:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 37:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 38:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 39:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=0;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 40:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 41:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 42:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 43:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 44:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 45:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 46:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 47:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 48:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 49:
 begin
    //Izquierda
    A7<=0;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 50:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 51:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 52:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 53:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 54:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 55:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 56:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 57:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1; 
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 58:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 59:
begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
end
 60:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 61:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 62:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 63:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 64:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 65:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 66:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 67:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 68:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 69:
 begin
    //Izquierda
    A7<=1;
    B7<=0;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 70:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 71:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 72:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 73:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 74:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 75:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 76:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 77:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 78:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 79:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=0;
    E7<=0;
    F7<=0;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 80:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 81:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 82:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 83:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;
 end
 84:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 85:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 86:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 87:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;   
 end
 88:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 89:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1; 
 end
 90:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
 91:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 92:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=0;
    D8<=1;
    E8<=1;
    F8<=0;
    G8<=1;
 end
 93:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=0;
    G8<=1;   
 end
 94:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=0;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 95:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 96:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=0;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 97:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=0;
    E8<=0;
    F8<=0;
    G8<=0;
 end
 98:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=1;
 end
 99:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=0;
    F7<=1;
    G7<=1;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=0;
    F8<=1;
    G8<=1;
 end
 default:
 begin
    //Izquierda
    A7<=1;
    B7<=1;
    C7<=1;
    D7<=1;
    E7<=1;
    F7<=1;
    G7<=0;
    //Derecha
    A8<=1;
    B8<=1;
    C8<=1;
    D8<=1;
    E8<=1;
    F8<=1;
    G8<=0;
 end
endcase
end
endmodule
