module Controlador_SEG(
    input [5:0] SEG,
    input CLK,
    input ALARM,
    //Digito Izquierda
    output reg A5,
    output reg B5,
    output reg C5,
    output reg D5,
    output reg E5,
    output reg F5,
    output reg G5,
    output reg DP5,
    //Digito Derecho
    output reg A6,
    output reg B6,
    output reg C6,
    output reg D6,
    output reg E6,
    output reg F6,
    output reg G6,
    output reg DP6
);
initial begin
    //Izquierda
    A5=0;
    B5=0;
    C5=0;
    D5=0;
    E5=0;
    F5=0;
    G5=0;
    DP5=0;
    //Derecha
    A6=0;
    B6=0;
    C6=0;
    D6=0;
    E6=0;
    F6=0;
    G6=0;
    DP6=1;
end

    reg[5:0] numero;

always @(posedge CLK)
begin
    if(ALARM)
    begin
        numero<=0;
    end
    else
    begin
        numero<=SEG;
    end
 case(numero)
 0:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 1:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 2:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 3:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;
 end
 4:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 5:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 6:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 7:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 8:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 9:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 10:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 11:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 12:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 13:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;
 end
 14:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 15:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 16:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 17:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 18:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 19:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=0;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 20:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 21:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 22:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 23:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;
 end
 24:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;  
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 25:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;  
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 26:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;  
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 27:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;  
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;   
 end
 28:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1;  
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 29:
 begin
     
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=0;
    D5<=1;
    E5<=1;
    F5<=0;
    G5<=1; 
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1; 
 end
 30:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 31:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 32:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 33:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;   
 end
 34:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 35:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 36:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 37:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 38:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 39:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=0;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 40:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 41:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 42:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 43:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;
 end
 44:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 45:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 46:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 47:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 48:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 49:
 begin
    //Izquierda
    A5<=0;
    B5<=1;
    C5<=1;
    D5<=0;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 50:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
 51:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 52:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=0;
    D6<=1;
    E6<=1;
    F6<=0;
    G6<=1;
 end
 53:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=0;
    G6<=1;
 end
 54:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=0;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 55:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
 end
 56:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=0;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 57:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1; 
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=0;
    E6<=0;
    F6<=0;
    G6<=0;
 end
 58:
 begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=1;
 end
 59:
begin
    //Izquierda
    A5<=1;
    B5<=0;
    C5<=1;
    D5<=1;
    E5<=0;
    F5<=1;
    G5<=1;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=0;
    F6<=1;
    G6<=1;
end
 default:
 begin
    //Izquierda
    A5<=1;
    B5<=1;
    C5<=1;
    D5<=1;
    E5<=1;
    F5<=1;
    G5<=0;
    //Derecha
    A6<=1;
    B6<=1;
    C6<=1;
    D6<=1;
    E6<=1;
    F6<=1;
    G6<=0;
 end
endcase
end
endmodule
