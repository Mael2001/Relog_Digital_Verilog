module Controlador_HORA(
    input [5:0] HORA,
    input CLK,
    input [5:0] AHORA,
    input ALARM,
    //Digito Izquierda
    output reg A1,
    output reg B1,
    output reg C1,
    output reg D1,
    output reg E1,
    output reg F1,
    output reg G1,
    output reg DP1,
    //Digito Derecho
    output reg A2,
    output reg B2,
    output reg C2,
    output reg D2,
    output reg E2,
    output reg F2,
    output reg G2,
    output reg DP2
);
initial begin
    //Izquierda
    A1=0;
    B1=0;
    C1=0;
    D1=0;
    E1=0;
    F1=0;
    G1=0;
    DP1=0;
    //Derecha
    A2=0;
    B2=0;
    C2=0;
    D2=0;
    E2=0;
    F2=0;
    G2=0;
    DP2=1;
end

    reg[5:0] numero;

always @(posedge CLK)
begin
    if(ALARM)
    begin
        numero<=AHORA;
    end
    else
    begin
        numero<=HORA;
    end
 case(numero)
 0:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=0;
 end
 1:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=0;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=0;
    G2<=0;
 end
 2:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=0;
    D2<=1;
    E2<=1;
    F2<=0;
    G2<=1;
 end
 3:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=0;
    G2<=1;
 end
 4:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=0;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 5:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=0;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 6:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=0;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=1;
 end
 7:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=0;
    G2<=0;
 end
 8:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=1;
 end
 9:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 10:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=0;
 end
 11:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=0;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=0;
    G2<=0;
 end
 12:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=0;
    D2<=1;
    E2<=1;
    F2<=0;
    G2<=1;
 end
 13:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=0;
    G2<=1;
 end
 14:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=0;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 15:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=0;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 16:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=0;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=1;
 end
 17:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=0;
    G2<=0;
 end
 18:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=1;
 end
 19:
 begin
    //Izquierda
    A1<=0;
    B1<=1;
    C1<=1;
    D1<=0;
    E1<=0;
    F1<=0;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=1;
    G2<=1;
 end
 20:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=0;
    D1<=1;
    E1<=1;
    F1<=0;
    G1<=1;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=0;
 end
 21:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=0;
    D1<=1;
    E1<=1;
    F1<=0;
    G1<=1;
    //Derecha
    A2<=0;
    B2<=1;
    C2<=1;
    D2<=0;
    E2<=0;
    F2<=0;
    G2<=0;
 end
 22:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=0;
    D1<=1;
    E1<=1;
    F1<=0;
    G1<=1;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=0;
    D2<=1;
    E2<=1;
    F2<=0;
    G2<=1;
 end
 23:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=0;
    D1<=1;
    E1<=1;
    F1<=0;
    G1<=1;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=0;
    F2<=0;
    G2<=1;
 end
 default:
 begin
    //Izquierda
    A1<=1;
    B1<=1;
    C1<=1;
    D1<=1;
    E1<=1;
    F1<=1;
    G1<=0;
    //Derecha
    A2<=1;
    B2<=1;
    C2<=1;
    D2<=1;
    E2<=1;
    F2<=1;
    G2<=0;
 end
endcase
end
endmodule
